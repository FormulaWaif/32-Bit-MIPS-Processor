----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:37:26 04/19/2024 
-- Design Name: 
-- Module Name:    Decoder - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Decoder is
    port (
        i: in std_logic_vector (4 downto 0); --input
		  write_ena: in std_logic; --enable of the decoder  
        o: out std_logic_vector (31 downto 0) --output
    );
end Decoder;

architecture rtl of Decoder is

begin
    o <= (OTHERS=>'Z') WHEN write_ena ='0' ELSE
    "00000000000000000000000000000001" WHEN i= "00000" ELSE
    "00000000000000000000000000000010" WHEN i= "00001" ELSE
    "00000000000000000000000000000100" WHEN i= "00010" ELSE
    "00000000000000000000000000001000" WHEN i= "00011" ELSE
    "00000000000000000000000000010000" WHEN i= "00100" ELSE
    "00000000000000000000000000100000" WHEN i= "00101" ELSE
    "00000000000000000000000001000000" WHEN i= "00110" ELSE
    "00000000000000000000000010000000" WHEN i= "00111" ELSE
    "00000000000000000000000100000000" WHEN i= "01000" ELSE
    "00000000000000000000001000000000" WHEN i= "01001" ELSE
    "00000000000000000000010000000000" WHEN i= "01010" ELSE
    "00000000000000000000100000000000" WHEN i= "01011" ELSE
    "00000000000000000001000000000000" WHEN i= "01100" ELSE
    "00000000000000000010000000000000" WHEN i= "01101" ELSE
    "00000000000000000100000000000000" WHEN i= "01110" ELSE
    "00000000000000001000000000000000" WHEN i= "01111" ELSE
    "00000000000000010000000000000000" WHEN i= "10000" ELSE
    "00000000000000100000000000000000" WHEN i= "10001" ELSE
    "00000000000001000000000000000000" WHEN i= "10010" ELSE
    "00000000000010000000000000000000" WHEN i= "10011" ELSE
    "00000000000100000000000000000000" WHEN i= "10100" ELSE
    "00000000001000000000000000000000" WHEN i= "10101" ELSE
    "00000000010000000000000000000000" WHEN i= "10110" ELSE
    "00000000100000000000000000000000" WHEN i= "10111" ELSE
    "00000001000000000000000000000000" WHEN i= "11000" ELSE
    "00000010000000000000000000000000" WHEN i= "11001" ELSE
    "00000100000000000000000000000000" WHEN i= "11010" ELSE
    "00001000000000000000000000000000" WHEN i= "11011" ELSE
    "00010000000000000000000000000000" WHEN i= "11100" ELSE
    "00100000000000000000000000000000" WHEN i= "11101" ELSE
    "01000000000000000000000000000000" WHEN i= "11110" ELSE
    "10000000000000000000000000000000" WHEN i= "11111" ELSE
    (OTHERS=>'Z');
end architecture;
